// This is our sequence

class seq1 extends uvm_sequence #(our_seq_item);
`uvm_object_utils(seq1)

function new(string name="seq1");
	super.new(name);
endfunction : new

//tasks


//

endclass : seq1