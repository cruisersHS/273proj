
module ebtb (
	input clk,
	input reset,
	input k,
	input [7:0] eb,
	output [9:0] tb,
	output reg disparity
);







endmodule : ebtb