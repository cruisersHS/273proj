//This is an empty sequencer


