//mimsg

class mimsg;
	reg [7:0] data;
endclass: mimsg
