
module crc32 (
	input clk,
	input reset,
	input [7:0] crc_in,
	input crc_in_valid,
	output [31:0] crc_out
);









endmodule : crc32